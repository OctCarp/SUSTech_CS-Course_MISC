`timescale 1ns / 1ps

module a2t4_dc (x, y);
    input[4: 0] x;
    output y;
    wire[3: 0]d10, d32;
    wire y0, y1, y2, y3, y4;
    
    d74139 dc10(0, x[1: 0], d10);
    d74139 dc32(0, x[3: 2], d32);
    
    and(y0, d10[3], d10[2], ~d10[1], d10[0], d32[3], d32[2], d32[1], ~d32[0], ~x[4]);
    and(y1, d10[3], ~d10[2], d10[1], d10[0], d32[3], d32[2], d32[1], ~d32[0], ~x[4]);
    and(y2, d10[3], d10[2], d10[1], ~d10[0], d32[3], d32[2], ~d32[1], d32[0], ~x[4]);
    and(y3, d10[3], d10[2], d10[1], ~d10[0], d32[3], ~d32[2], d32[1], d32[0], ~x[4]);
    and(y4, d10[3], d10[2], d10[1], ~d10[0], d32[3], d32[2], d32[1], ~d32[0], x[4]);
    
    or(y, y0, y1, y2, y3, y4);
endmodule
